library verilog;
use verilog.vl_types.all;
entity lab6fsm_vlg_vec_tst is
end lab6fsm_vlg_vec_tst;
