library verilog;
use verilog.vl_types.all;
entity ALUProblem3_vlg_vec_tst is
end ALUProblem3_vlg_vec_tst;
