library verilog;
use verilog.vl_types.all;
entity ALUProblem2_vlg_vec_tst is
end ALUProblem2_vlg_vec_tst;
