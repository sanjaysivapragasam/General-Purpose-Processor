library verilog;
use verilog.vl_types.all;
entity ssegmodified_vlg_vec_tst is
end ssegmodified_vlg_vec_tst;
