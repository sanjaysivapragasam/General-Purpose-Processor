library verilog;
use verilog.vl_types.all;
entity ALUproblem1_vlg_vec_tst is
end ALUproblem1_vlg_vec_tst;
